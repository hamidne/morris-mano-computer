module ALU(Data, AC, AND, DR, ADD, DR, INPR, INPT, COM, SHL, E, SHR);
	input [15:0] AC, DR;
	input [7:0] INPR;
	input  AND, ADD, DR, INPR, INPT, COM, SHL, E, SHR ;
	