module FGO_FlipFlop();

endmodule