module IEN_FlipFlop();

endmodule